library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity microcode_rom is

end microcode_rom;

architecture Behavioral of microcode_rom is

begin


end Behavioral;
