
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity control_unit is
--  Port ( );
end control_unit;

architecture Behavioral of control_unit is

begin


end Behavioral;
